`define     V48_ON                         16'hb201 
`define     V48_ENABLE                     16'hb20c 
`define     K1_ON                          16'hb202 
`define     K1_ENABLE                      16'hb20d 
`define     AUX_FAN_CTL                    16'hb203 
`define     AUX_0_CTL                      16'hb204 
`define     AUX_1_CTL                      16'hb205 
`define     AUX_2_CTL                      16'hb206 
`define     AUX_3_CTL                      16'hb207 
`define     RESET                          16'hb208 
`define     CTR_CTL                        16'hb209 
`define     GEN_FREQ_CTR_MUX               16'hb227 
`define     V0_LO                          16'hb20a 
`define     V0_HI                          16'hb20b 
`define     I1_LO                          16'hb210 
`define     I1_HI                          16'hb211 
`define     I2_LO                          16'hb212 
`define     I2_HI                          16'hb213 
`define     MAIN_BLOWER_LO                 16'hb21e 
`define     MAIN_BLOWER_HI                 16'hb21f 
`define     GEN_FREQ_CTR_LO                16'hb228 
`define     GEN_FREQ_CTR_MID               16'hb226 
`define     GEN_FREQ_CTR_HI                16'hb229 
`define     BC_TACH0_CTR_LO                16'hb22d 
`define     BC_TACH0_CTR_HI                16'hb22e 
`define     BC_TACH1_CTR_LO                16'hb22f 
`define     BC_TACH1_CTR_HI                16'hb230 
`define     BC_TACH_CTL                    16'hb231 
`define     ID_REV                         16'hb22a 
`define     MAINT_MON                      16'hb22b 
`define     LOCK_OUT_STATE                 16'hb22c 
`define     B_CNTRL_BC_48VDC               16'hb301 
`define     B_DC90_48V_Enable              16'hb30c 
`define     B_CNTRL_BC_48VDC_DC90          16'hb304 
`define     DC90_STATE                     16'hb32e 
`define     STATE_48V                      16'hb32b 
`define     STATE_BC_FAN                   16'hb310 
`define     B_SMC_CNTRL_BC_SWITCHED_AC     16'hb305 
`define     SMC_MON_BC_AC_ON               16'hb32a 
`define     SMC_CNTRL_JAG_SWITCHED_AC      16'hb302 
`define     SMC_MON_PDU_K1                 16'hb303 
`define     SMC_CNTRL_JAG_48VDC_ON         16'hb306 
`define     SMC_MON_PDU_JAG_48V_GOOD       16'hb311 
`define     SMC_MON_PDU_JAG_48V_LVL_ON     16'hb32c 
`define     SMC_MON_PDU_JAG_THERMAL_FAULT  16'hb30a 
